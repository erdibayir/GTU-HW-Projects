library verilog;
use verilog.vl_types.all;
entity mips32_tb is
    port(
        testout         : out    vl_logic
    );
end mips32_tb;
