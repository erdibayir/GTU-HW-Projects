module sub_32_bit(i1,i2,out);
input [31:0] i1,i2;
output [31:0] out;
wire a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,a32;
wire cout;
wire b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15,b16,b17,b18,b19,b20,b21,b22,b23,b24,b25,b26,b27,b28,b29,b30,b31,b32;

xor(a1,i1[0],1);
xor(a2,i1[1],1);
xor(a3,i1[2],1);
xor(a4,i1[3],1);
xor(a5,i1[4],1);
xor(a6,i1[5],1);
xor(a7,i1[6],1);
xor(a8,i1[7],1);
xor(a9,i1[8],1);
xor(a10,i1[9],1);
xor(a11,i1[10],1);
xor(a12,i1[11],1);
xor(a13,i1[12],1);
xor(a14,i1[13],1);
xor(a15,i1[14],1);
xor(a16,i1[15],1);
xor(a17,i1[16],1);
xor(a18,i1[17],1);
xor(a19,i1[18],1);
xor(a20,i1[19],1);
xor(a21,i1[20],1);
xor(a22,i1[21],1);
xor(a23,i1[22],1);
xor(a24,i1[23],1);
xor(a25,i1[24],1);
xor(a26,i1[25],1);
xor(a27,i1[26],1);
xor(a28,i1[27],1);
xor(a29,i1[28],1);
xor(a30,i1[29],1);
xor(a31,i1[30],1);
xor(a32,i1[31],1);


full_adder f1(a1,i2[0],1'b0,b1,cout);
full_adder f2(a2,i2[1],cout,b2,cout1);
full_adder f3(a3,i2[2],cout1,b3,cout2);
full_adder f4(a4,i2[3],cout2,b4,cout3);
full_adder f5(a5,i2[4],cout3,b5,cout4);
full_adder f6(a6,i2[5],cout4,b6,cout5);
full_adder f7(a7,i2[6],cout5,b7,cout6);
full_adder f8(a8,i2[7],cout6,b8,cout7);
full_adder f9(a9,i2[8],cout7,b9,cout8);
full_adder f10(a10,i2[9],cout8,b10,cout9);
full_adder f11(a11,i2[10],cout9,b11,cout10);
full_adder f12(a12,i2[11],cout10,b12,cout11);
full_adder f13(a13,i2[12],cout11,b13,cout12);
full_adder f14(a14,i2[13],cout12,b14,cout13);
full_adder f15(a15,i2[14],cout13,b15,cout14);
full_adder f16(a16,i2[15],cout14,b16,cout15);
full_adder f17(a17,i2[16],cout15,b17,cout16);
full_adder f18(a18,i2[17],cout16,b18,cout17);
full_adder f19(a19,i2[18],cout17,b19,cout18);
full_adder f20(a20,i2[19],cout18,b20,cout19);
full_adder f21(a21,i2[20],cout19,b21,cout20);
full_adder f22(a22,i2[21],cout20,b22,cout21);
full_adder f23(a23,i2[22],cout21,b23,cout22);
full_adder f24(a24,i2[23],cout22,b24,cout23);
full_adder f25(a25,i2[24],cout23,b25,cout24);
full_adder f26(a26,i2[25],cout24,b26,cout25);
full_adder f27(a27,i2[26],cout25,b27,cout26);
full_adder f28(a28,i2[27],cout26,b28,cout27);
full_adder f29(a29,i2[28],cout27,b29,cout28);
full_adder f30(a30,i2[29],cout28,b30,cout29);
full_adder f31(a31,i2[30],cout29,b31,cout30);
full_adder f32(a32,i2[31],cout30,b32,cout31);

not(out[0],b1);
not(out[1],b2);
not(out[2],b3);
not(out[3],b4);
not(out[4],b5);
not(out[5],b6);
not(out[6],b7);
not(out[7],b8);
not(out[8],b9);
not(out[9],b10);
not(out[10],b11);
not(out[11],b12);
not(out[12],b13);
not(out[13],b14);
not(out[14],b15);
not(out[15],b16);
not(out[16],b17);
not(out[17],b18);
not(out[18],b19);
not(out[19],b20);
not(out[20],b21);
not(out[21],b22);
not(out[22],b23);
not(out[23],b24);
not(out[24],b25);
not(out[25],b26);
not(out[26],b27);
not(out[27],b28);
not(out[28],b29);
not(out[29],b30);
not(out[30],b31);
not(out[31],b32);

endmodule