module or_32_bit(i1,i2,out);

input [31:0] i1,i2;
output [31:0] out;

or x1(out[0],i1[0],i2[0]);
or x2(out[1],i1[1],i2[1]);
or x3(out[2],i1[2],i2[2]);
or x4(out[3],i1[3],i2[3]);
or x5(out[4],i1[4],i2[4]);
or x6(out[5],i1[5],i2[5]);
or x7(out[6],i1[6],i2[6]);
or x8(out[7],i1[7],i2[7]);
or x9(out[8],i1[8],i2[8]);
or x10(out[9],i1[9],i2[9]);
or x11(out[10],i1[10],i2[10]);
or x12(out[11],i1[11],i2[11]);
or x13(out[12],i1[12],i2[12]);
or x14(out[13],i1[13],i2[13]);
or x15(out[14],i1[14],i2[14]);
or x16(out[15],i1[15],i2[15]);
or x17(out[16],i1[16],i2[16]);
or x18(out[17],i1[17],i2[17]);
or x19(out[18],i1[18],i2[18]);
or x20(out[19],i1[19],i2[19]);
or x21(out[20],i1[20],i2[20]);
or x22(out[21],i1[21],i2[21]);
or x23(out[22],i1[22],i2[22]);
or x24(out[23],i1[23],i2[23]);
or x25(out[24],i1[24],i2[24]);
or x26(out[25],i1[25],i2[25]);
or x27(out[26],i1[26],i2[26]);
or x28(out[27],i1[27],i2[27]);
or x29(out[28],i1[28],i2[28]);
or x30(out[29],i1[29],i2[29]);
or x31(out[30],i1[30],i2[30]);
or x32(out[31],i1[31],i2[31]);

endmodule